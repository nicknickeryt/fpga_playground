`timescale 1ns / 1ps
module 7seg(
input  [3:0] a,
output [3:0] y
    );

y[0] = 1'b1;

endmodule